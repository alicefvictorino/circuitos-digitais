ENTITY decodificador_portas_logicas IS
port(
A1, A2, A3, A4: in bit;
S0, S1, S2, S3, S4, S5, S6: out bit);
END;

ARCHITECTURE behav OF decodificador_portas_logicas IS
BEGIN
S0 <= (NOT A1 AND NOT A2 AND A3 AND NOT A4) OR (A1 AND NOT A2 AND NOT A3 AND NOT A4);
S1 <= (A1 AND NOT A2 AND A3 AND NOT A4) OR (NOT A1 AND A2 AND A3 AND NOT A4);
S2 <= NOT A1 AND A2 AND NOT A3 AND NOT A4;
S3 <= (A1 AND NOT A2 AND NOT A3 AND NOT A4) OR (NOT A1 AND NOT A2 AND A3 AND NOT A4)
OR (A1 AND A2 AND A3 AND NOT A4);
S4 <= (A1 AND A2 AND NOT A4) OR (A1 AND NOT A2 AND NOT A3) OR (NOT A2 AND A3 AND NOT
A4);
S5 <= (A1 AND A2 AND NOT A4) OR (A2 AND NOT A3 AND NOT A4) OR (A1 AND NOT A3 AND NOT
A4);
S6 <= (A1 AND A2 AND A3 AND NOT A4) OR (NOT A2 AND NOT A3 AND NOT A4);
END;
